module control_unit(
    
)